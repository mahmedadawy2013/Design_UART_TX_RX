library verilog;
use verilog.vl_types.all;
entity UART_TX_tb is
end UART_TX_tb;
